`timescale 1ns/1ps

module RCA_8bitTestbench;



endmodule


