`timescale 1ns/1ps

module Mem_To_Reg_Selector(
    input [31:0] ,
    input [31:0] ,
    input [31:0] prog_count,
    output reg [31:0] data_write,

)